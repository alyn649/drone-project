library verilog;
use verilog.vl_types.all;
entity drone_vlg_vec_tst is
end drone_vlg_vec_tst;
